library ieee;
use ieee.std_logic_1164.all;

entity tristate_dr is
	port
	(
		d_in  : in std_logic_vector(7 downto 0);
		en    : in std_logic;
		d_out : out std_logic_vector(7 downto 0);
		rst   : in std_logic
	);
end tristate_dr;

architecture behavior of tristate_dr is
	signal local_signal : std_logic;
begin

	tristate_driver : process (d_in, en)
		variable local_variable_tristate : std_logic := '0';
	begin
		if en = '1' then
			d_out <= d_in;
		else
			-- array can be created simply by using vector
			d_out <= "ZZZZZZZZ";
		end if;
	end process tristate_driver;

	p_rst : process (rst)
	begin
		if rst = '1' then
			local_signal <= '0';
		end if;
	end process;

end behavior;